module Shifter( dataA, dataB, Signal, dataOut, reset );
input reset ;
input [31:0] dataA ;
input [4:0] dataB ;
input [5:0] Signal ;
output [31:0] dataOut ;

wire [31:0] temp0, temp1, temp2, temp3, temp ;

parameter SRL = 6'b000010;

    Mux221 U_mux221_11(.sel(dataB[0]), .a(dataA[0]), .b(dataA[1]), .y(temp0[0]) );
    Mux221 U_mux221_12(.sel(dataB[0]), .a(dataA[1]), .b(dataA[2]), .y(temp0[1]) );
    Mux221 U_mux221_13(.sel(dataB[0]), .a(dataA[2]), .b(dataA[3]), .y(temp0[2]) );
    Mux221 U_mux221_14(.sel(dataB[0]), .a(dataA[3]), .b(dataA[4]), .y(temp0[3]) );
    Mux221 U_mux221_15(.sel(dataB[0]), .a(dataA[4]), .b(dataA[5]), .y(temp0[4]) );
    Mux221 U_mux221_16(.sel(dataB[0]), .a(dataA[5]), .b(dataA[6]), .y(temp0[5]) );
    Mux221 U_mux221_17(.sel(dataB[0]), .a(dataA[6]), .b(dataA[7]), .y(temp0[6]) );
    Mux221 U_mux221_18(.sel(dataB[0]), .a(dataA[7]), .b(dataA[8]), .y(temp0[7]) );
    Mux221 U_mux221_19(.sel(dataB[0]), .a(dataA[8]), .b(dataA[9]), .y(temp0[8]) );
    Mux221 U_mux221_10(.sel(dataB[0]), .a(dataA[9]), .b(dataA[10]), .y(temp0[9]) );
    Mux221 U_mux221_111(.sel(dataB[0]), .a(dataA[10]), .b(dataA[11]), .y(temp0[10]) );
    Mux221 U_mux221_112(.sel(dataB[0]), .a(dataA[11]), .b(dataA[12]), .y(temp0[11]) );
    Mux221 U_mux221_113(.sel(dataB[0]), .a(dataA[12]), .b(dataA[13]), .y(temp0[12]) );
    Mux221 U_mux221_114(.sel(dataB[0]), .a(dataA[13]), .b(dataA[14]), .y(temp0[13]) );
    Mux221 U_mux221_115(.sel(dataB[0]), .a(dataA[14]), .b(dataA[15]), .y(temp0[14]) );
    Mux221 U_mux221_116(.sel(dataB[0]), .a(dataA[15]), .b(dataA[16]), .y(temp0[15]) );
    Mux221 U_mux221_117(.sel(dataB[0]), .a(dataA[16]), .b(dataA[17]), .y(temp0[16]) );
    Mux221 U_mux221_118(.sel(dataB[0]), .a(dataA[17]), .b(dataA[18]), .y(temp0[17]) );
    Mux221 U_mux221_119(.sel(dataB[0]), .a(dataA[18]), .b(dataA[19]), .y(temp0[18]) );
    Mux221 U_mux221_120(.sel(dataB[0]), .a(dataA[19]), .b(dataA[20]), .y(temp0[19]) );
    Mux221 U_mux221_121(.sel(dataB[0]), .a(dataA[20]), .b(dataA[21]), .y(temp0[20]) );
    Mux221 U_mux221_122(.sel(dataB[0]), .a(dataA[21]), .b(dataA[22]), .y(temp0[21]) );
    Mux221 U_mux221_123(.sel(dataB[0]), .a(dataA[22]), .b(dataA[23]), .y(temp0[22]) );
    Mux221 U_mux221_124(.sel(dataB[0]), .a(dataA[23]), .b(dataA[24]), .y(temp0[23]) );
    Mux221 U_mux221_125(.sel(dataB[0]), .a(dataA[24]), .b(dataA[25]), .y(temp0[24]) );
    Mux221 U_mux221_126(.sel(dataB[0]), .a(dataA[25]), .b(dataA[26]), .y(temp0[25]) );
    Mux221 U_mux221_127(.sel(dataB[0]), .a(dataA[26]), .b(dataA[27]), .y(temp0[26]) );
    Mux221 U_mux221_128(.sel(dataB[0]), .a(dataA[27]), .b(dataA[28]), .y(temp0[27]) );
    Mux221 U_mux221_129(.sel(dataB[0]), .a(dataA[28]), .b(dataA[29]), .y(temp0[28]) );
    Mux221 U_mux221_130(.sel(dataB[0]), .a(dataA[29]), .b(dataA[30]), .y(temp0[29]) );
    Mux221 U_mux221_131(.sel(dataB[0]), .a(dataA[30]), .b(dataA[31]), .y(temp0[30]) );
    Mux221 U_mux221_132(.sel(dataB[0]), .a(dataA[31]), .b(1'b0), .y(temp0[31]) );
    
    Mux221 U_mux221_21(.sel(dataB[1]), .a(temp0[0]), .b(temp0[2]), .y(temp1[0]) );
    Mux221 U_mux221_22(.sel(dataB[1]), .a(temp0[1]), .b(temp0[3]), .y(temp1[1]) );
    Mux221 U_mux221_23(.sel(dataB[1]), .a(temp0[2]), .b(temp0[4]), .y(temp1[2]) );
    Mux221 U_mux221_24(.sel(dataB[1]), .a(temp0[3]), .b(temp0[5]), .y(temp1[3]) );
    Mux221 U_mux221_25(.sel(dataB[1]), .a(temp0[4]), .b(temp0[6]), .y(temp1[4]) );
    Mux221 U_mux221_26(.sel(dataB[1]), .a(temp0[5]), .b(temp0[7]), .y(temp1[5]) );
    Mux221 U_mux221_27(.sel(dataB[1]), .a(temp0[6]), .b(temp0[8]), .y(temp1[6]) );
    Mux221 U_mux221_28(.sel(dataB[1]), .a(temp0[7]), .b(temp0[9]), .y(temp1[7]) );
    Mux221 U_mux221_29(.sel(dataB[1]), .a(temp0[8]), .b(temp0[10]), .y(temp1[8]) );
    Mux221 U_mux221_20(.sel(dataB[1]), .a(temp0[9]), .b(temp0[11]), .y(temp1[9]) );
    Mux221 U_mux221_211(.sel(dataB[1]), .a(temp0[10]), .b(temp0[12]), .y(temp1[10]) );
    Mux221 U_mux221_212(.sel(dataB[1]), .a(temp0[11]), .b(temp0[13]), .y(temp1[11]) );
    Mux221 U_mux221_213(.sel(dataB[1]), .a(temp0[12]), .b(temp0[14]), .y(temp1[12]) );
    Mux221 U_mux221_214(.sel(dataB[1]), .a(temp0[13]), .b(temp0[15]), .y(temp1[13]) );
    Mux221 U_mux221_215(.sel(dataB[1]), .a(temp0[14]), .b(temp0[16]), .y(temp1[14]) );
    Mux221 U_mux221_216(.sel(dataB[1]), .a(temp0[15]), .b(temp0[17]), .y(temp1[15]) );
    Mux221 U_mux221_217(.sel(dataB[1]), .a(temp0[16]), .b(temp0[18]), .y(temp1[16]) );
    Mux221 U_mux221_218(.sel(dataB[1]), .a(temp0[17]), .b(temp0[19]), .y(temp1[17]) );
    Mux221 U_mux221_219(.sel(dataB[1]), .a(temp0[18]), .b(temp0[20]), .y(temp1[18]) );
    Mux221 U_mux221_220(.sel(dataB[1]), .a(temp0[19]), .b(temp0[21]), .y(temp1[19]) );
    Mux221 U_mux221_221(.sel(dataB[1]), .a(temp0[20]), .b(temp0[22]), .y(temp1[20]) );
    Mux221 U_mux221_222(.sel(dataB[1]), .a(temp0[21]), .b(temp0[23]), .y(temp1[21]) );
    Mux221 U_mux221_223(.sel(dataB[1]), .a(temp0[22]), .b(temp0[24]), .y(temp1[22]) );
    Mux221 U_mux221_224(.sel(dataB[1]), .a(temp0[23]), .b(temp0[25]), .y(temp1[23]) );
    Mux221 U_mux221_225(.sel(dataB[1]), .a(temp0[24]), .b(temp0[26]), .y(temp1[24]) );
    Mux221 U_mux221_226(.sel(dataB[1]), .a(temp0[25]), .b(temp0[27]), .y(temp1[25]) );
    Mux221 U_mux221_227(.sel(dataB[1]), .a(temp0[26]), .b(temp0[28]), .y(temp1[26]) );
    Mux221 U_mux221_228(.sel(dataB[1]), .a(temp0[27]), .b(temp0[29]), .y(temp1[27]) );
    Mux221 U_mux221_229(.sel(dataB[1]), .a(temp0[28]), .b(temp0[30]), .y(temp1[28]) );
    Mux221 U_mux221_230(.sel(dataB[1]), .a(temp0[29]), .b(temp0[31]), .y(temp1[29]) );
    Mux221 U_mux221_231(.sel(dataB[1]), .a(temp0[30]), .b(1'b0), .y(temp1[30]) );
    Mux221 U_mux221_232(.sel(dataB[1]), .a(temp0[31]), .b(1'b0), .y(temp1[31]) );
  
    Mux221 U_mux221_31(.sel(dataB[2]), .a(temp1[0]), .b(temp1[4]), .y(temp2[0]) );
    Mux221 U_mux221_32(.sel(dataB[2]), .a(temp1[1]), .b(temp1[5]), .y(temp2[1]) );
    Mux221 U_mux221_33(.sel(dataB[2]), .a(temp1[2]), .b(temp1[6]), .y(temp2[2]) );
    Mux221 U_mux221_34(.sel(dataB[2]), .a(temp1[3]), .b(temp1[7]), .y(temp2[3]) );
    Mux221 U_mux221_35(.sel(dataB[2]), .a(temp1[4]), .b(temp1[8]), .y(temp2[4]) );
    Mux221 U_mux221_36(.sel(dataB[2]), .a(temp1[5]), .b(temp1[9]), .y(temp2[5]) );
    Mux221 U_mux221_37(.sel(dataB[2]), .a(temp1[6]), .b(temp1[10]), .y(temp2[6]) );
    Mux221 U_mux221_38(.sel(dataB[2]), .a(temp1[7]), .b(temp1[11]), .y(temp2[7]) );
    Mux221 U_mux221_39(.sel(dataB[2]), .a(temp1[8]), .b(temp1[12]), .y(temp2[8]) );
    Mux221 U_mux221_30(.sel(dataB[2]), .a(temp1[9]), .b(temp1[13]), .y(temp2[9]) );
    Mux221 U_mux221_311(.sel(dataB[2]), .a(temp1[10]), .b(temp1[14]), .y(temp2[10]) );
    Mux221 U_mux221_312(.sel(dataB[2]), .a(temp1[11]), .b(temp1[15]), .y(temp2[11]) );
    Mux221 U_mux221_313(.sel(dataB[2]), .a(temp1[12]), .b(temp1[16]), .y(temp2[12]) );
    Mux221 U_mux221_314(.sel(dataB[2]), .a(temp1[13]), .b(temp1[17]), .y(temp2[13]) );
    Mux221 U_mux221_315(.sel(dataB[2]), .a(temp1[14]), .b(temp1[18]), .y(temp2[14]) );
    Mux221 U_mux221_316(.sel(dataB[2]), .a(temp1[15]), .b(temp1[19]), .y(temp2[15]) );
    Mux221 U_mux221_317(.sel(dataB[2]), .a(temp1[16]), .b(temp1[20]), .y(temp2[16]) );
    Mux221 U_mux221_318(.sel(dataB[2]), .a(temp1[17]), .b(temp1[21]), .y(temp2[17]) );
    Mux221 U_mux221_319(.sel(dataB[2]), .a(temp1[18]), .b(temp1[22]), .y(temp2[18]) );
    Mux221 U_mux221_320(.sel(dataB[2]), .a(temp1[19]), .b(temp1[23]), .y(temp2[19]) );
    Mux221 U_mux221_321(.sel(dataB[2]), .a(temp1[20]), .b(temp1[24]), .y(temp2[20]) );
    Mux221 U_mux221_322(.sel(dataB[2]), .a(temp1[21]), .b(temp1[25]), .y(temp2[21]) );
    Mux221 U_mux221_323(.sel(dataB[2]), .a(temp1[22]), .b(temp1[26]), .y(temp2[22]) );
    Mux221 U_mux221_324(.sel(dataB[2]), .a(temp1[23]), .b(temp1[27]), .y(temp2[23]) );
    Mux221 U_mux221_325(.sel(dataB[2]), .a(temp1[24]), .b(temp1[28]), .y(temp2[24]) );
    Mux221 U_mux221_326(.sel(dataB[2]), .a(temp1[25]), .b(temp1[29]), .y(temp2[25]) );
    Mux221 U_mux221_327(.sel(dataB[2]), .a(temp1[26]), .b(temp1[30]), .y(temp2[26]) );
    Mux221 U_mux221_328(.sel(dataB[2]), .a(temp1[27]), .b(temp1[31]), .y(temp2[27]) );
    Mux221 U_mux221_329(.sel(dataB[2]), .a(temp1[28]), .b(1'b0), .y(temp2[28]) );
    Mux221 U_mux221_330(.sel(dataB[2]), .a(temp1[29]), .b(1'b0), .y(temp2[29]) );
    Mux221 U_mux221_331(.sel(dataB[2]), .a(temp1[30]), .b(1'b0), .y(temp2[30]) );
    Mux221 U_mux221_332(.sel(dataB[2]), .a(temp1[31]), .b(1'b0), .y(temp2[31]) );
    
    Mux221 U_mux221_41(.sel(dataB[3]), .a(temp2[0]), .b(temp2[8]), .y(temp3[0]) );
    Mux221 U_mux221_42(.sel(dataB[3]), .a(temp2[1]), .b(temp2[9]), .y(temp3[1]) );
    Mux221 U_mux221_43(.sel(dataB[3]), .a(temp2[2]), .b(temp2[10]), .y(temp3[2]) );
    Mux221 U_mux221_44(.sel(dataB[3]), .a(temp2[3]), .b(temp2[11]), .y(temp3[3]) );
    Mux221 U_mux221_45(.sel(dataB[3]), .a(temp2[4]), .b(temp2[12]), .y(temp3[4]) );
    Mux221 U_mux221_46(.sel(dataB[3]), .a(temp2[5]), .b(temp2[13]), .y(temp3[5]) );
    Mux221 U_mux221_47(.sel(dataB[3]), .a(temp2[6]), .b(temp2[14]), .y(temp3[6]) );
    Mux221 U_mux221_48(.sel(dataB[3]), .a(temp2[7]), .b(temp2[15]), .y(temp3[7]) );
    Mux221 U_mux221_49(.sel(dataB[3]), .a(temp2[8]), .b(temp2[16]), .y(temp3[8]) );
    Mux221 U_mux221_40(.sel(dataB[3]), .a(temp2[9]), .b(temp2[17]), .y(temp3[9]) );
    Mux221 U_mux221_411(.sel(dataB[3]), .a(temp2[10]), .b(temp2[18]), .y(temp3[10]) );
    Mux221 U_mux221_412(.sel(dataB[3]), .a(temp2[11]), .b(temp2[19]), .y(temp3[11]) );
    Mux221 U_mux221_413(.sel(dataB[3]), .a(temp2[12]), .b(temp2[20]), .y(temp3[12]) );
    Mux221 U_mux221_414(.sel(dataB[3]), .a(temp2[13]), .b(temp2[21]), .y(temp3[13]) );
    Mux221 U_mux221_415(.sel(dataB[3]), .a(temp2[14]), .b(temp2[22]), .y(temp3[14]) );
    Mux221 U_mux221_416(.sel(dataB[3]), .a(temp2[15]), .b(temp2[23]), .y(temp3[15]) );
    Mux221 U_mux221_417(.sel(dataB[3]), .a(temp2[16]), .b(temp2[24]), .y(temp3[16]) );
    Mux221 U_mux221_418(.sel(dataB[3]), .a(temp2[17]), .b(temp2[25]), .y(temp3[17]) );
    Mux221 U_mux221_419(.sel(dataB[3]), .a(temp2[18]), .b(temp2[26]), .y(temp3[18]) );
    Mux221 U_mux221_420(.sel(dataB[3]), .a(temp2[19]), .b(temp2[27]), .y(temp3[19]) );
    Mux221 U_mux221_421(.sel(dataB[3]), .a(temp2[20]), .b(temp2[28]), .y(temp3[20]) );
    Mux221 U_mux221_422(.sel(dataB[3]), .a(temp2[21]), .b(temp2[29]), .y(temp3[21]) );
    Mux221 U_mux221_423(.sel(dataB[3]), .a(temp2[22]), .b(temp2[30]), .y(temp3[22]) );
    Mux221 U_mux221_424(.sel(dataB[3]), .a(temp2[23]), .b(temp2[31]), .y(temp3[23]) );
    Mux221 U_mux221_425(.sel(dataB[3]), .a(temp2[24]), .b(1'b0), .y(temp3[24]) );
    Mux221 U_mux221_426(.sel(dataB[3]), .a(temp2[25]), .b(1'b0), .y(temp3[25]) );
    Mux221 U_mux221_427(.sel(dataB[3]), .a(temp2[26]), .b(1'b0), .y(temp3[26]) );
    Mux221 U_mux221_428(.sel(dataB[3]), .a(temp2[27]), .b(1'b0), .y(temp3[27]) );
    Mux221 U_mux221_429(.sel(dataB[3]), .a(temp2[28]), .b(1'b0), .y(temp3[28]) );
    Mux221 U_mux221_430(.sel(dataB[3]), .a(temp2[29]), .b(1'b0), .y(temp3[29]) );
    Mux221 U_mux221_431(.sel(dataB[3]), .a(temp2[30]), .b(1'b0), .y(temp3[30]) );
    Mux221 U_mux221_432(.sel(dataB[3]), .a(temp2[31]), .b(1'b0), .y(temp3[31]) );
  
    Mux221 U_mux221_51(.sel(dataB[4]), .a(temp3[0]), .b(temp3[16]), .y(temp[0]) );
    Mux221 U_mux221_52(.sel(dataB[4]), .a(temp3[1]), .b(temp3[17]), .y(temp[1]) );
    Mux221 U_mux221_53(.sel(dataB[4]), .a(temp3[2]), .b(temp3[18]), .y(temp[2]) );
    Mux221 U_mux221_54(.sel(dataB[4]), .a(temp3[3]), .b(temp3[19]), .y(temp[3]) );
    Mux221 U_mux221_55(.sel(dataB[4]), .a(temp3[4]), .b(temp3[20]), .y(temp[4]) );
    Mux221 U_mux221_56(.sel(dataB[4]), .a(temp3[5]), .b(temp3[21]), .y(temp[5]) );
    Mux221 U_mux221_57(.sel(dataB[4]), .a(temp3[6]), .b(temp3[22]), .y(temp[6]) );
    Mux221 U_mux221_58(.sel(dataB[4]), .a(temp3[7]), .b(temp3[23]), .y(temp[7]) );
    Mux221 U_mux221_59(.sel(dataB[4]), .a(temp3[8]), .b(temp3[24]), .y(temp[8]) );
    Mux221 U_mux221_50(.sel(dataB[4]), .a(temp3[9]), .b(temp3[25]), .y(temp[9]) );
    Mux221 U_mux221_511(.sel(dataB[4]), .a(temp3[10]), .b(temp3[26]), .y(temp[10]) );
    Mux221 U_mux221_512(.sel(dataB[4]), .a(temp3[11]), .b(temp3[27]), .y(temp[11]) );
    Mux221 U_mux221_513(.sel(dataB[4]), .a(temp3[12]), .b(temp3[28]), .y(temp[12]) );
    Mux221 U_mux221_514(.sel(dataB[4]), .a(temp3[13]), .b(temp3[29]), .y(temp[13]) );
    Mux221 U_mux221_515(.sel(dataB[4]), .a(temp3[14]), .b(temp3[30]), .y(temp[14]) );
    Mux221 U_mux221_516(.sel(dataB[4]), .a(temp3[15]), .b(temp3[31]), .y(temp[15]) );
    Mux221 U_mux221_517(.sel(dataB[4]), .a(temp3[16]), .b(1'b0), .y(temp[16]) );
    Mux221 U_mux221_518(.sel(dataB[4]), .a(temp3[17]), .b(1'b0), .y(temp[17]) );
    Mux221 U_mux221_519(.sel(dataB[4]), .a(temp3[18]), .b(1'b0), .y(temp[18]) );
    Mux221 U_mux221_520(.sel(dataB[4]), .a(temp3[19]), .b(1'b0), .y(temp[19]) );
    Mux221 U_mux221_521(.sel(dataB[4]), .a(temp3[20]), .b(1'b0), .y(temp[20]) );
    Mux221 U_mux221_522(.sel(dataB[4]), .a(temp3[21]), .b(1'b0), .y(temp[21]) );
    Mux221 U_mux221_523(.sel(dataB[4]), .a(temp3[22]), .b(1'b0), .y(temp[22]) );
    Mux221 U_mux221_524(.sel(dataB[4]), .a(temp3[23]), .b(1'b0), .y(temp[23]) );
    Mux221 U_mux221_525(.sel(dataB[4]), .a(temp3[24]), .b(1'b0), .y(temp[24]) );
    Mux221 U_mux221_526(.sel(dataB[4]), .a(temp3[25]), .b(1'b0), .y(temp[25]) );
    Mux221 U_mux221_527(.sel(dataB[4]), .a(temp3[26]), .b(1'b0), .y(temp[26]) );
    Mux221 U_mux221_528(.sel(dataB[4]), .a(temp3[27]), .b(1'b0), .y(temp[27]) );
    Mux221 U_mux221_529(.sel(dataB[4]), .a(temp3[28]), .b(1'b0), .y(temp[28]) );
    Mux221 U_mux221_530(.sel(dataB[4]), .a(temp3[29]), .b(1'b0), .y(temp[29]) );
    Mux221 U_mux221_531(.sel(dataB[4]), .a(temp3[30]), .b(1'b0), .y(temp[30]) );
    Mux221 U_mux221_532(.sel(dataB[4]), .a(temp3[31]), .b(1'b0), .y(temp[31]) );
  
      
  
assign dataOut = reset ? 32'b0 : (Signal== SRL) ? temp : dataOut ;

endmodule

	
